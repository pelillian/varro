module pin_out (
p_out, p_in); 

output p_out;
input p_in; 

assign p_out = p_in; 

endmodule
